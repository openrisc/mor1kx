/* ****************************************************************************
  This Source Code Form is subject to the terms of the
  Open Hardware Description License, v. 1.0. If a copy
  of the OHDL was not distributed with this file, You
  can obtain one at http://juliusbaxter.net/ohdl/ohdl.txt

  Description: mor1kx branch control

  Muxes between branches from decode stage and branches generated by
  exceptions.
  Copyright (C) 2012 - 2013 Authors

   Author(s): Julius Baxter <juliusbaxter@gmail.com>
              Stefan Kristiansson <stefan.kristiansson@saunalahti.fi>

***************************************************************************** */

`include "mor1kx-defines.v"

module mor1kx_ctrl_branch_cappuccino
  #(
    parameter OPTION_OPERAND_WIDTH = 32
    )
   (
    input 			      clk,
    input 			      rst,

    // Inputs from decode stage
    input 			      decode_branch_i,
    input [OPTION_OPERAND_WIDTH-1:0]  decode_branch_target_i,

    input 			      ctrl_branch_exception_i,
    input [OPTION_OPERAND_WIDTH-1:0]  ctrl_branch_except_pc_i,

    input 			      ctrl_except_syscall_i,

    output 			      ctrl_branch_occur_o,
    output [OPTION_OPERAND_WIDTH-1:0] ctrl_branch_target_o
    );



   // Exceptions take precedence
   assign ctrl_branch_occur_o = ctrl_branch_exception_i |
				/* we have to prevent branches when we have
				 * syscall exception in control stage
				 * TODO: check if there are other exceptions
				 * that need this too */
				!ctrl_except_syscall_i & decode_branch_i;


   assign ctrl_branch_target_o = ctrl_branch_exception_i ?
				 ctrl_branch_except_pc_i :
				 decode_branch_target_i;

endmodule // mor1kx_ctrl_branch_cappuccino
