/*
 mor1kx processor top level
 */

`include "mor1kx-defines.v"

module mor1kx
  (/*AUTOARG*/
   // Outputs
   iwbm_adr_o, iwbm_stb_o, iwbm_cyc_o, iwbm_sel_o, iwbm_we_o,
   iwbm_cti_o, iwbm_bte_o, iwbm_dat_o, dwbm_adr_o, dwbm_stb_o,
   dwbm_cyc_o, dwbm_sel_o, dwbm_we_o, dwbm_cti_o, dwbm_bte_o,
   dwbm_dat_o, du_dat_o, du_ack_o, du_stall_o,
   // Inputs
   clk, rst, iwbm_err_i, iwbm_ack_i, iwbm_dat_i, iwbm_rty_i,
   dwbm_err_i, dwbm_ack_i, dwbm_dat_i, dwbm_rty_i, irq_i, du_addr_i,
   du_stb_i, du_dat_i, du_we_i, du_stall_i
   );

   parameter OPTION_OPERAND_WIDTH = 32;

   parameter OPTION_CPU0 = "FOURSTAGE";

   parameter FEATURE_DATACACHE = "NONE";
   parameter OPTION_DCACHE_BLOCK_WIDTH = 5;
   parameter OPTION_DCACHE_SET_WIDTH = 9;
   parameter OPTION_DCACHE_WAYS = 2;
   parameter OPTION_DCACHE_LIMIT_WIDTH = 32;
   parameter FEATURE_DMMU = "NONE";
   parameter FEATURE_INSTRUCTIONCACHE = "NONE";
   parameter OPTION_ICACHE_BLOCK_WIDTH = 5;
   parameter OPTION_ICACHE_SET_WIDTH = 9;
   parameter OPTION_ICACHE_WAYS = 2;
   parameter OPTION_ICACHE_LIMIT_WIDTH = 32;
   parameter FEATURE_IMMU = "NONE";
   parameter FEATURE_PIC = "ENABLED";
   parameter FEATURE_TIMER = "ENABLED";
   parameter FEATURE_DEBUGUNIT = "NONE";
   parameter FEATURE_PERFCOUNTERS = "NONE";
   parameter FEATURE_MAC = "NONE";

   parameter FEATURE_SYSCALL = "ENABLED";
   parameter FEATURE_TRAP = "ENABLED";
   parameter FEATURE_RANGE = "ENABLED";

   parameter OPTION_PIC_TRIGGER = "EDGE";

   parameter OPTION_RF_ADDR_WIDTH = 5;
   parameter OPTION_RF_WORDS = 32;

   parameter OPTION_RESET_PC = {{(OPTION_OPERAND_WIDTH-13){1'b0}},
				`OR1K_RESET_VECTOR,8'd0};

   parameter FEATURE_MULTIPLIER = "THREESTAGE";
   parameter FEATURE_DIVIDER = "SERIAL";

   parameter FEATURE_ADDC = "NONE";
   parameter FEATURE_SRA = "ENABLED";
   parameter FEATURE_ROR = "NONE";
   parameter FEATURE_EXT = "NONE";
   parameter FEATURE_CMOV = "NONE";
   parameter FEATURE_FFL1 = "ENABLED";
   
   parameter FEATURE_CUST1 = "NONE";
   parameter FEATURE_CUST2 = "NONE";
   parameter FEATURE_CUST3 = "NONE";
   parameter FEATURE_CUST4 = "NONE";
   parameter FEATURE_CUST5 = "NONE";
   parameter FEATURE_CUST6 = "NONE";
   parameter FEATURE_CUST7 = "NONE";
   parameter FEATURE_CUST8 = "NONE";
   
   parameter OPTION_SHIFTER = "BARREL";

   parameter BUS_IF_TYPE = "WISHBONE32";
   
   input clk, rst;
   
   output [31:0] iwbm_adr_o;
   output 	 iwbm_stb_o;
   output 	 iwbm_cyc_o;
   output [3:0]  iwbm_sel_o;
   output 	 iwbm_we_o;
   output [2:0]  iwbm_cti_o;
   output [1:0]  iwbm_bte_o;
   output [31:0] iwbm_dat_o;
   input 	 iwbm_err_i;
   input 	 iwbm_ack_i;
   input [31:0]  iwbm_dat_i;
   input 	 iwbm_rty_i;

   output [31:0] dwbm_adr_o;
   output 	 dwbm_stb_o;
   output 	 dwbm_cyc_o;
   output [3:0]  dwbm_sel_o;
   output 	 dwbm_we_o;
   output [2:0]  dwbm_cti_o;
   output [1:0]  dwbm_bte_o;
   output [31:0] dwbm_dat_o;
   input 	 dwbm_err_i;
   input 	 dwbm_ack_i;
   input [31:0]  dwbm_dat_i;
   input 	 dwbm_rty_i;

   input [31:0]  irq_i;

   // Debug interface
   input [15:0]  du_addr_i;
   input 	 du_stb_i;
   input [OPTION_OPERAND_WIDTH-1:0] du_dat_i;
   input 			    du_we_i;
   output [OPTION_OPERAND_WIDTH-1:0] du_dat_o;
   output 			     du_ack_o;
   // Stall control from debug interface
   input 			     du_stall_i;
   output 			     du_stall_o;
   

   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire [OPTION_OPERAND_WIDTH-1:0] dbus_adr_o;	// From mor1kx_cpu of mor1kx_cpu.v
   wire [3:0]		dbus_bsel_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire [OPTION_OPERAND_WIDTH-1:0] dbus_dat_o;	// From mor1kx_cpu of mor1kx_cpu.v
   wire			dbus_req_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire			dbus_we_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire			dc_ack_i;		// From dbus_bridge of mor1kx_bus_if_wb32.v
   wire [OPTION_OPERAND_WIDTH-1:0] dc_dat_i;	// From dbus_bridge of mor1kx_bus_if_wb32.v
   wire			dc_err_i;		// From dbus_bridge of mor1kx_bus_if_wb32.v
   wire [OPTION_OPERAND_WIDTH-1:0] ibus_adr_o;	// From mor1kx_cpu of mor1kx_cpu.v
   wire			ibus_req_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire			ic_ack_i;		// From ibus_bridge of mor1kx_bus_if_wb32.v
   wire [`OR1K_INSN_WIDTH-1:0] ic_dat_i;	// From ibus_bridge of mor1kx_bus_if_wb32.v
   wire			ic_err_i;		// From ibus_bridge of mor1kx_bus_if_wb32.v
   wire			spr_bus_ack_dc_i;	// From mor1kx_dcache of mor1kx_dcache.v
   wire			spr_bus_ack_ic_i;	// From mor1kx_icache of mor1kx_icache.v
   wire [15:0]		spr_bus_addr_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire [OPTION_OPERAND_WIDTH-1:0] spr_bus_dat_dc_i;// From mor1kx_dcache of mor1kx_dcache.v
   wire [OPTION_OPERAND_WIDTH-1:0] spr_bus_dat_ic_i;// From mor1kx_icache of mor1kx_icache.v
   wire [OPTION_OPERAND_WIDTH-1:0] spr_bus_dat_o;// From mor1kx_cpu of mor1kx_cpu.v
   wire			spr_bus_stb_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire			spr_bus_we_o;		// From mor1kx_cpu of mor1kx_cpu.v
   wire [15:0]		spr_sr_o;		// From mor1kx_cpu of mor1kx_cpu.v
   // End of automatics

   wire 			   ibus_ack_i;
   wire [OPTION_OPERAND_WIDTH-1:0] ibus_dat_i;
   wire 			   ibus_err_i;
   wire [OPTION_OPERAND_WIDTH-1:0] ic_adr_o;
   wire 			   ic_req_o;

   wire 			   dbus_ack_i;
   wire [OPTION_OPERAND_WIDTH-1:0] dbus_dat_i;
   wire 			   dbus_err_i;
   wire [OPTION_OPERAND_WIDTH-1:0] dc_adr_o;
   wire 			   dc_req_o;
   wire 			   dc_we_o;
   wire [OPTION_OPERAND_WIDTH-1:0] dc_dat_o;
   wire [3:0] 			   dc_bsel_o;

   generate
      if (BUS_IF_TYPE=="WISHBONE32") begin : bus_gen

	 /* mor1kx_bus_if_wb32 AUTO_TEMPLATE (
	  .cpu_err_o			(ic_err_i),
	  .cpu_ack_o			(ic_ack_i),
	  .cpu_dat_o			(ic_dat_i[`OR1K_INSN_WIDTH-1:0]),
	  .wbm_adr_o			(iwbm_adr_o),
	  .wbm_stb_o			(iwbm_stb_o),
	  .wbm_cyc_o			(iwbm_cyc_o),
	  .wbm_sel_o			(iwbm_sel_o),
	  .wbm_we_o			(iwbm_we_o),
	  .wbm_cti_o			(iwbm_cti_o),
	  .wbm_bte_o			(iwbm_bte_o),
	  .wbm_dat_o			(iwbm_dat_o),
	  // Inputs
	  .cpu_adr_i			(ic_adr_o),
	  .cpu_dat_i			(0),
	  .cpu_req_i			(ic_req_o),
	  .cpu_we_i			(0),
	  .cpu_bsel_i			(4'b1111),
	  .wbm_err_i			(iwbm_err_i),
	  .wbm_ack_i			(iwbm_ack_i),
	  .wbm_dat_i			(iwbm_dat_i),
	  .wbm_rty_i			(iwbm_rty_i),
	  ); */
	 
	 mor1kx_bus_if_wb32 
//		      #(.BUS_IF_TYPE("CLASSIC"))
		      #(.BUS_IF_TYPE("B3_READ_BURSTING"))
	 ibus_bridge
		      (/*AUTOINST*/
		       // Outputs
		       .cpu_err_o	(ic_err_i),		 // Templated
		       .cpu_ack_o	(ic_ack_i),		 // Templated
		       .cpu_dat_o	(ic_dat_i[`OR1K_INSN_WIDTH-1:0]), // Templated
		       .wbm_adr_o	(iwbm_adr_o),		 // Templated
		       .wbm_stb_o	(iwbm_stb_o),		 // Templated
		       .wbm_cyc_o	(iwbm_cyc_o),		 // Templated
		       .wbm_sel_o	(iwbm_sel_o),		 // Templated
		       .wbm_we_o	(iwbm_we_o),		 // Templated
		       .wbm_cti_o	(iwbm_cti_o),		 // Templated
		       .wbm_bte_o	(iwbm_bte_o),		 // Templated
		       .wbm_dat_o	(iwbm_dat_o),		 // Templated
		       // Inputs
		       .clk		(clk),
		       .rst		(rst),
		       .cpu_adr_i	(ic_adr_o),		 // Templated
		       .cpu_dat_i	(0),			 // Templated
		       .cpu_req_i	(ic_req_o),		 // Templated
		       .cpu_bsel_i	(4'b1111),		 // Templated
		       .cpu_we_i	(0),			 // Templated
		       .wbm_err_i	(iwbm_err_i),		 // Templated
		       .wbm_ack_i	(iwbm_ack_i),		 // Templated
		       .wbm_dat_i	(iwbm_dat_i),		 // Templated
		       .wbm_rty_i	(iwbm_rty_i));		 // Templated
	 
	 /* mor1kx_bus_if_wb32 AUTO_TEMPLATE (
	  .cpu_err_o			(dc_err_i),
	  .cpu_ack_o			(dc_ack_i),
	  .cpu_dat_o			(dc_dat_i[OPTION_OPERAND_WIDTH-1:0]),
	  .wbm_adr_o			(dwbm_adr_o),
	  .wbm_stb_o			(dwbm_stb_o),
	  .wbm_cyc_o			(dwbm_cyc_o),
	  .wbm_sel_o			(dwbm_sel_o),
	  .wbm_we_o			(dwbm_we_o),
	  .wbm_cti_o			(dwbm_cti_o),
	  .wbm_bte_o			(dwbm_bte_o),
	  .wbm_dat_o			(dwbm_dat_o),
	  // Inputs
	  .cpu_adr_i			(dc_adr_o[31:0]),
	  .cpu_dat_i			(dc_dat_o),
	  .cpu_req_i			(dc_req_o),
	  .cpu_we_i			(dc_we_o),
	  .cpu_bsel_i			(dc_bsel_o),
	  .wbm_err_i			(dwbm_err_i),
	  .wbm_ack_i			(dwbm_ack_i),
	  .wbm_dat_i			(dwbm_dat_i),
	  .wbm_rty_i			(dwbm_rty_i),
	  ); */

	 mor1kx_bus_if_wb32
	   #(.BUS_IF_TYPE("CLASSIC"))
	 dbus_bridge
	   (/*AUTOINST*/
	    // Outputs
	    .cpu_err_o			(dc_err_i),		 // Templated
	    .cpu_ack_o			(dc_ack_i),		 // Templated
	    .cpu_dat_o			(dc_dat_i[OPTION_OPERAND_WIDTH-1:0]), // Templated
	    .wbm_adr_o			(dwbm_adr_o),		 // Templated
	    .wbm_stb_o			(dwbm_stb_o),		 // Templated
	    .wbm_cyc_o			(dwbm_cyc_o),		 // Templated
	    .wbm_sel_o			(dwbm_sel_o),		 // Templated
	    .wbm_we_o			(dwbm_we_o),		 // Templated
	    .wbm_cti_o			(dwbm_cti_o),		 // Templated
	    .wbm_bte_o			(dwbm_bte_o),		 // Templated
	    .wbm_dat_o			(dwbm_dat_o),		 // Templated
	    // Inputs
	    .clk			(clk),
	    .rst			(rst),
	    .cpu_adr_i			(dc_adr_o[31:0]),	 // Templated
	    .cpu_dat_i			(dc_dat_o),		 // Templated
	    .cpu_req_i			(dc_req_o),		 // Templated
	    .cpu_bsel_i			(dc_bsel_o),		 // Templated
	    .cpu_we_i			(dc_we_o),		 // Templated
	    .wbm_err_i			(dwbm_err_i),		 // Templated
	    .wbm_ack_i			(dwbm_ack_i),		 // Templated
	    .wbm_dat_i			(dwbm_dat_i),		 // Templated
	    .wbm_rty_i			(dwbm_rty_i));		 // Templated
	 
      end // if (BUS_IF_TYPE=="WISHBONE32")
      else
	begin
	   initial begin
	      $display("Error: BUS_IF_TYPE not correct");
	      $finish();
	   end
	end // else: !if(BUS_IF_TYPE=="WISHBONE32")
   endgenerate

   generate
      if (FEATURE_INSTRUCTIONCACHE!="NONE") begin : icache_gen

   /* mor1kx_icache AUTO_TEMPLATE (
	    // Outputs
	    .cpu_err_o			(ibus_err_i),
	    .cpu_ack_o			(ibus_ack_i),
	    .cpu_dat_o			(ibus_dat_i[31:0]),
	    .spr_bus_dat_o		(spr_bus_dat_ic_i[OPTION_OPERAND_WIDTH-1:0]),
	    .spr_bus_ack_o		(spr_bus_ack_ic_i),
	    // Inputs
	    .ic_enable			(spr_sr_o[`OR1K_SPR_SR_ICE]),
	    .cpu_adr_i			(ibus_adr_o[31:0]),
	    .cpu_req_i			(ibus_req_o),
	    .spr_bus_addr_i		(spr_bus_addr_o[15:0]),
	    .spr_bus_we_i		(spr_bus_we_o),
	    .spr_bus_stb_i		(spr_bus_stb_o),
	    .spr_bus_dat_i		(spr_bus_dat_o[OPTION_OPERAND_WIDTH-1:0]),
    );*/

   mor1kx_icache
     #(
       .OPTION_ICACHE_BLOCK_WIDTH(OPTION_ICACHE_BLOCK_WIDTH),
       .OPTION_ICACHE_SET_WIDTH(OPTION_ICACHE_SET_WIDTH),
       .OPTION_ICACHE_WAYS(OPTION_ICACHE_WAYS),
       .OPTION_ICACHE_LIMIT_WIDTH(OPTION_ICACHE_LIMIT_WIDTH)
       )
   mor1kx_icache
	   (/*AUTOINST*/
	    // Outputs
	    .cpu_err_o			(ibus_err_i),		 // Templated
	    .cpu_ack_o			(ibus_ack_i),		 // Templated
	    .cpu_dat_o			(ibus_dat_i[31:0]),	 // Templated
	    .ic_adr_o			(ic_adr_o[31:0]),
	    .ic_req_o			(ic_req_o),
	    .spr_bus_dat_o		(spr_bus_dat_ic_i[OPTION_OPERAND_WIDTH-1:0]), // Templated
	    .spr_bus_ack_o		(spr_bus_ack_ic_i),	 // Templated
	    // Inputs
	    .clk			(clk),
	    .rst			(rst),
	    .ic_enable			(spr_sr_o[`OR1K_SPR_SR_ICE]), // Templated
	    .cpu_adr_i			(ibus_adr_o[31:0]),	 // Templated
	    .cpu_req_i			(ibus_req_o),		 // Templated
	    .ic_err_i			(ic_err_i),
	    .ic_ack_i			(ic_ack_i),
	    .ic_dat_i			(ic_dat_i[31:0]),
	    .spr_bus_addr_i		(spr_bus_addr_o[15:0]),	 // Templated
	    .spr_bus_we_i		(spr_bus_we_o),		 // Templated
	    .spr_bus_stb_i		(spr_bus_stb_o),	 // Templated
	    .spr_bus_dat_i		(spr_bus_dat_o[OPTION_OPERAND_WIDTH-1:0])); // Templated
      end
      else
	begin
	   assign ibus_ack_i = ic_ack_i;
	   assign ibus_dat_i = ic_dat_i;
	   assign ibus_err_i = ic_err_i;
	   assign ic_adr_o = ibus_adr_o;
	   assign ic_req_o = ibus_req_o;
	end
   endgenerate

   generate
      if (FEATURE_DATACACHE!="NONE") begin : dcache_gen

   /* mor1kx_dcache AUTO_TEMPLATE (
	    // Outputs
	    .cpu_err_o			(dbus_err_i),
	    .cpu_ack_o			(dbus_ack_i),
	    .cpu_dat_o			(dbus_dat_i[31:0]),
	    .spr_bus_dat_o		(spr_bus_dat_dc_i[OPTION_OPERAND_WIDTH-1:0]),
	    .spr_bus_ack_o		(spr_bus_ack_dc_i),
	    // Inputs
	    .dc_enable			(spr_sr_o[`OR1K_SPR_SR_DCE]),
	    .cpu_dat_i			(dbus_dat_o[31:0]),
	    .cpu_adr_i			(dbus_adr_o[31:0]),
	    .cpu_req_i			(dbus_req_o),
	    .cpu_we_i			(dbus_we_o),
	    .cpu_bsel_i			(dbus_bsel_o[3:0]),
	    .spr_bus_addr_i		(spr_bus_addr_o[15:0]),
	    .spr_bus_we_i		(spr_bus_we_o),
	    .spr_bus_stb_i		(spr_bus_stb_o),
	    .spr_bus_dat_i		(spr_bus_dat_o[OPTION_OPERAND_WIDTH-1:0]),
    );*/

   mor1kx_dcache
     #(
       .OPTION_DCACHE_BLOCK_WIDTH(OPTION_DCACHE_BLOCK_WIDTH),
       .OPTION_DCACHE_SET_WIDTH(OPTION_DCACHE_SET_WIDTH),
       .OPTION_DCACHE_WAYS(OPTION_DCACHE_WAYS),
       .OPTION_DCACHE_LIMIT_WIDTH(OPTION_DCACHE_LIMIT_WIDTH)
       )
   mor1kx_dcache
	   (/*AUTOINST*/
	    // Outputs
	    .cpu_err_o			(dbus_err_i),		 // Templated
	    .cpu_ack_o			(dbus_ack_i),		 // Templated
	    .cpu_dat_o			(dbus_dat_i[31:0]),	 // Templated
	    .dc_dat_o			(dc_dat_o[31:0]),
	    .dc_adr_o			(dc_adr_o[31:0]),
	    .dc_req_o			(dc_req_o),
	    .dc_we_o			(dc_we_o),
	    .dc_bsel_o			(dc_bsel_o[3:0]),
	    .spr_bus_dat_o		(spr_bus_dat_dc_i[OPTION_OPERAND_WIDTH-1:0]), // Templated
	    .spr_bus_ack_o		(spr_bus_ack_dc_i),	 // Templated
	    // Inputs
	    .clk			(clk),
	    .rst			(rst),
	    .dc_enable			(spr_sr_o[`OR1K_SPR_SR_DCE]), // Templated
	    .cpu_dat_i			(dbus_dat_o[31:0]),	 // Templated
	    .cpu_adr_i			(dbus_adr_o[31:0]),	 // Templated
	    .cpu_req_i			(dbus_req_o),		 // Templated
	    .cpu_we_i			(dbus_we_o),		 // Templated
	    .cpu_bsel_i			(dbus_bsel_o[3:0]),	 // Templated
	    .dc_err_i			(dc_err_i),
	    .dc_ack_i			(dc_ack_i),
	    .dc_dat_i			(dc_dat_i[31:0]),
	    .spr_bus_addr_i		(spr_bus_addr_o[15:0]),	 // Templated
	    .spr_bus_we_i		(spr_bus_we_o),		 // Templated
	    .spr_bus_stb_i		(spr_bus_stb_o),	 // Templated
	    .spr_bus_dat_i		(spr_bus_dat_o[OPTION_OPERAND_WIDTH-1:0])); // Templated
      end
      else
	begin
	   assign dbus_ack_i = dc_ack_i;
	   assign dbus_dat_i = dc_dat_i;
	   assign dbus_err_i = dc_err_i;
	   assign dc_adr_o = dbus_adr_o;
	   assign dc_req_o = dbus_req_o;
	   assign dc_we_o = dbus_we_o;
	   assign dc_dat_o = dbus_dat_o;
	   assign dc_bsel_o = dbus_bsel_o;
	end
   endgenerate

   /* mor1kx_cpu AUTO_TEMPLATE
    ( .spr_bus_dat_dc_i		(),
    .spr_bus_ack_dc_i		(),
    .spr_bus_dat_ic_i		(spr_bus_dat_ic_i),
    .spr_bus_ack_ic_i		(spr_bus_ack_ic_i),
    .spr_bus_dat_dmmu_i		(),
    .spr_bus_ack_dmmu_i		(),
    .spr_bus_dat_immu_i		(),
    .spr_bus_ack_immu_i		(),
    .spr_bus_dat_mac_i		(),
    .spr_bus_ack_mac_i		(),
    .spr_bus_dat_pmu_i		(),
    .spr_bus_ack_pmu_i		(),
    .spr_bus_dat_pcu_i		(),
    .spr_bus_ack_pcu_i		(),
    .spr_bus_dat_fpu_i		(),
    .spr_bus_ack_fpu_i		(),
    ); */
   mor1kx_cpu  
     	   #(
	     .OPTION_OPERAND_WIDTH(OPTION_OPERAND_WIDTH),
	     .OPTION_CPU(OPTION_CPU0),
	     .FEATURE_DATACACHE(FEATURE_DATACACHE),
	     .OPTION_DCACHE_BLOCK_WIDTH(OPTION_DCACHE_BLOCK_WIDTH),
	     .OPTION_DCACHE_SET_WIDTH(OPTION_DCACHE_SET_WIDTH),
	     .OPTION_DCACHE_WAYS(OPTION_DCACHE_WAYS),
	     .FEATURE_DMMU(FEATURE_DMMU),
	     .FEATURE_INSTRUCTIONCACHE(FEATURE_INSTRUCTIONCACHE),
	     .OPTION_ICACHE_BLOCK_WIDTH(OPTION_ICACHE_BLOCK_WIDTH),
	     .OPTION_ICACHE_SET_WIDTH(OPTION_ICACHE_SET_WIDTH),
	     .OPTION_ICACHE_WAYS(OPTION_ICACHE_WAYS),
	     .FEATURE_IMMU(FEATURE_IMMU),
	     .FEATURE_PIC(FEATURE_PIC),
	     .FEATURE_TIMER(FEATURE_TIMER),
	     .FEATURE_DEBUGUNIT(FEATURE_DEBUGUNIT),
	     .FEATURE_PERFCOUNTERS(FEATURE_PERFCOUNTERS),
	     .FEATURE_MAC(FEATURE_MAC),
	     .FEATURE_SYSCALL(FEATURE_SYSCALL),
	     .FEATURE_TRAP(FEATURE_TRAP),
	     .FEATURE_RANGE(FEATURE_RANGE),
	     .OPTION_PIC_TRIGGER(OPTION_PIC_TRIGGER),
	     .OPTION_RF_ADDR_WIDTH(OPTION_RF_ADDR_WIDTH),
	     .OPTION_RF_WORDS(OPTION_RF_WORDS),
	     .OPTION_RESET_PC(OPTION_RESET_PC),
	     .FEATURE_MULTIPLIER(FEATURE_MULTIPLIER),
	     .FEATURE_DIVIDER(FEATURE_DIVIDER),
	     .FEATURE_ADDC(FEATURE_ADDC),
	     .FEATURE_SRA(FEATURE_SRA),
	     .FEATURE_ROR(FEATURE_ROR),
	     .FEATURE_EXT(FEATURE_EXT),
	     .FEATURE_CMOV(FEATURE_CMOV),
	     .FEATURE_FFL1(FEATURE_FFL1),
	     .FEATURE_CUST1(FEATURE_CUST1),
	     .FEATURE_CUST2(FEATURE_CUST2),
	     .FEATURE_CUST3(FEATURE_CUST3),
	     .FEATURE_CUST4(FEATURE_CUST4),
	     .FEATURE_CUST5(FEATURE_CUST5),
	     .FEATURE_CUST6(FEATURE_CUST6),
	     .FEATURE_CUST7(FEATURE_CUST7),
	     .FEATURE_CUST8(FEATURE_CUST8),
	     .OPTION_SHIFTER(OPTION_SHIFTER)
	     )
   mor1kx_cpu
     (/*AUTOINST*/
      // Outputs
      .ibus_adr_o			(ibus_adr_o[OPTION_OPERAND_WIDTH-1:0]),
      .ibus_req_o			(ibus_req_o),
      .dbus_adr_o			(dbus_adr_o[OPTION_OPERAND_WIDTH-1:0]),
      .dbus_dat_o			(dbus_dat_o[OPTION_OPERAND_WIDTH-1:0]),
      .dbus_req_o			(dbus_req_o),
      .dbus_bsel_o			(dbus_bsel_o[3:0]),
      .dbus_we_o			(dbus_we_o),
      .du_dat_o				(du_dat_o[OPTION_OPERAND_WIDTH-1:0]),
      .du_ack_o				(du_ack_o),
      .du_stall_o			(du_stall_o),
      .spr_bus_addr_o			(spr_bus_addr_o[15:0]),
      .spr_bus_we_o			(spr_bus_we_o),
      .spr_bus_stb_o			(spr_bus_stb_o),
      .spr_bus_dat_o			(spr_bus_dat_o[OPTION_OPERAND_WIDTH-1:0]),
      .spr_sr_o				(spr_sr_o[15:0]),
      // Inputs
      .clk				(clk),
      .rst				(rst),
      .ibus_err_i			(ibus_err_i),
      .ibus_ack_i			(ibus_ack_i),
      .ibus_dat_i			(ibus_dat_i[`OR1K_INSN_WIDTH-1:0]),
      .dbus_err_i			(dbus_err_i),
      .dbus_ack_i			(dbus_ack_i),
      .dbus_dat_i			(dbus_dat_i[OPTION_OPERAND_WIDTH-1:0]),
      .irq_i				(irq_i[31:0]),
      .du_addr_i			(du_addr_i[15:0]),
      .du_stb_i				(du_stb_i),
      .du_dat_i				(du_dat_i[OPTION_OPERAND_WIDTH-1:0]),
      .du_we_i				(du_we_i),
      .du_stall_i			(du_stall_i),
      .spr_bus_dat_dc_i			(),			 // Templated
      .spr_bus_ack_dc_i			(),			 // Templated
      .spr_bus_dat_ic_i			(spr_bus_dat_ic_i),	 // Templated
      .spr_bus_ack_ic_i			(spr_bus_ack_ic_i),	 // Templated
      .spr_bus_dat_dmmu_i		(),			 // Templated
      .spr_bus_ack_dmmu_i		(),			 // Templated
      .spr_bus_dat_immu_i		(),			 // Templated
      .spr_bus_ack_immu_i		(),			 // Templated
      .spr_bus_dat_mac_i		(),			 // Templated
      .spr_bus_ack_mac_i		(),			 // Templated
      .spr_bus_dat_pmu_i		(),			 // Templated
      .spr_bus_ack_pmu_i		(),			 // Templated
      .spr_bus_dat_pcu_i		(),			 // Templated
      .spr_bus_ack_pcu_i		(),			 // Templated
      .spr_bus_dat_fpu_i		(),			 // Templated
      .spr_bus_ack_fpu_i		());			 // Templated
   
endmodule // mor1kx
