/******************************************************************************
 This Source Code Form is subject to the terms of the
 Open Hardware Description License, v. 1.0. If a copy
 of the OHDL was not distributed with this file, You
 can obtain one at http://juliusbaxter.net/ohdl/ohdl.txt

 Description: Single port ram

 Copyright (C) 2012 Stefan Kristiansson <stefan.kristiansson@saunalahti.fi>

 ******************************************************************************/

module mor1kx_spram
  #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32
    )
   (
    input 		    clk,
    input [ADDR_WIDTH-1:0]  raddr,
    input [ADDR_WIDTH-1:0]  waddr,
    input 		    we,
    input [DATA_WIDTH-1:0]  din,
    output [DATA_WIDTH-1:0] dout
    );

   reg [DATA_WIDTH-1:0]     mem[(1<<ADDR_WIDTH)-1:0];
   reg [DATA_WIDTH-1:0]     rdata;
   reg [DATA_WIDTH-1:0]     din_r;

   reg 			    bypass;

   assign dout = bypass ? din_r : rdata;

   always @(posedge clk) begin
      if (we)
	mem[waddr] <= din;
      rdata <= mem[raddr];
   end

   always @(posedge clk)
     din_r <= din;

   always @(posedge clk)
     if (waddr == raddr && we)
       bypass <= 1;
     else
       bypass <= 0;

endmodule
